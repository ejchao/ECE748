package decode_in_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "src/decode_in_transaction.svh"
    `include "src/decode_in_coverage.svh"
    `include "src/decode_in_configuration.svh"
    `include "src/decode_in_sequence_base.svh"
    `include "src/decode_in_random_sequence.svh"
    `include "src/decode_in_monitor.svh"
    `include "src/decode_in_driver.svh"
    `include "src/decode_in_agent.svh"

endpackage