package decode_test_pkg;

    import uvmf_base_pkg::*;
    import uvmf_base_pkg_hdl::*;
    import uvm_pkg::*;
    import decode_in_pkg::*;
    import decode_out_pkg::*;
    `include "uvm_macros.svh"
    `include "src/test_top.svh"
    //`include "src/print_component.svh"

endpackage